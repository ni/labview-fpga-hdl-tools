-------------------------------------------------------------------------------
--
-- File: PkgLvFpgaConst.vhd
-- Original Project: Puma 1.5
-- Date: 24 Jan 2008
--
-------------------------------------------------------------------------------
-- (c) 2008 Copyright National Instruments Corporation
-- All Rights Reserved
-- National Instruments Internal Information
-------------------------------------------------------------------------------
--
-- Purpose:
--  This file will be generated by LV FPGA to set constants required for
--  Puma 1.5 compilation.
--
-------------------------------------------------------------------------------

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package PkgLvFpgaConst is

  -----------------------------------------------------------------------------
  -- LV FPGA generated constants
  -----------------------------------------------------------------------------

  constant kExpectedTbId   : std_logic_vector(31 downto 0) := X"10937AEC";
  constant kExpectDumbTb   : std_logic := '0';
  constant kEnableFamClockSync : std_logic := '1';
  constant kFamClockSrcSel  : std_logic := '1';
  constant kInsertBank0Mig  : boolean := false;
  constant kInsertBank1Mig  : boolean := false;
  constant kInsertHostMemoryBufferMig  : boolean := false;
  constant kInsertLowLatencyBufferMig  : boolean := false;
  constant kAuxMgtClipPresent  : boolean :=  false;
  constant kAuxDioDefaultVoltage : natural := 3300;
  constant kCfgSubsysId : std_logic_vector(15 downto 0) := X"7AEC";
  constant kDram2DPBaseAddress : natural := 16#20000#;
  
end PkgLvFpgaConst;

package body PkgLvFpgaConst is

  
end PkgLvFpgaConst;

