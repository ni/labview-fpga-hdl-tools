----------------------------------------------
-- IMPLEMENTATION NOT NEEDED FOR TESTING
----------------------------------------------