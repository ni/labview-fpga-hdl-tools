xIoModuleReady <= xIoModuleReady;
xIoModuleErrorCode <= xIoModuleErrorCode;
aDioOut <= aDioOut;
aDioIn <= aDioIn;
UserClkPort0 <= UserClkPort0;
aPort0PmaInit <= aPort0PmaInit;
aPort0ResetPb <= aPort0ResetPb;
uPort0AxiTxTData0 <= uPort0AxiTxTData0;
uPort0AxiTxTData1 <= uPort0AxiTxTData1;
uPort0AxiTxTData2 <= uPort0AxiTxTData2;
uPort0AxiTxTData3 <= uPort0AxiTxTData3;
uPort0AxiTxTKeep <= uPort0AxiTxTKeep;
uPort0AxiTxTLast <= uPort0AxiTxTLast;
uPort0AxiTxTValid <= uPort0AxiTxTValid;
uPort0AxiTxTReady <= uPort0AxiTxTReady;
uPort0AxiRxTData0 <= uPort0AxiRxTData0;
uPort0AxiRxTData1 <= uPort0AxiRxTData1;
uPort0AxiRxTData2 <= uPort0AxiRxTData2;
uPort0AxiRxTData3 <= uPort0AxiRxTData3;
uPort0AxiRxTKeep <= uPort0AxiRxTKeep;
uPort0AxiRxTLast <= uPort0AxiRxTLast;
uPort0AxiRxTValid <= uPort0AxiRxTValid;
uPort0AxiNfcTValid <= uPort0AxiNfcTValid;
uPort0AxiNfcTData <= uPort0AxiNfcTData;
uPort0AxiNfcTReady <= uPort0AxiNfcTReady;
uPort0HardError <= uPort0HardError;
uPort0SoftError <= uPort0SoftError;
uPort0LaneUp <= uPort0LaneUp;
uPort0ChannelUp <= uPort0ChannelUp;
uPort0SysResetOut <= uPort0SysResetOut;
uPort0MmcmNotLockOut <= uPort0MmcmNotLockOut;
uPort0CrcPassFail_n <= uPort0CrcPassFail_n;
uPort0CrcValid <= uPort0CrcValid;
iPort0LinkResetOut <= iPort0LinkResetOut;
sGtwiz0CtrlAxiAWAddr <= sGtwiz0CtrlAxiAWAddr;
sGtwiz0CtrlAxiAWValid <= sGtwiz0CtrlAxiAWValid;
sGtwiz0CtrlAxiAWReady <= sGtwiz0CtrlAxiAWReady;
sGtwiz0CtrlAxiWData <= sGtwiz0CtrlAxiWData;
sGtwiz0CtrlAxiWStrb <= sGtwiz0CtrlAxiWStrb;
sGtwiz0CtrlAxiWValid <= sGtwiz0CtrlAxiWValid;
sGtwiz0CtrlAxiWReady <= sGtwiz0CtrlAxiWReady;
sGtwiz0CtrlAxiBResp <= sGtwiz0CtrlAxiBResp;
sGtwiz0CtrlAxiBValid <= sGtwiz0CtrlAxiBValid;
sGtwiz0CtrlAxiBReady <= sGtwiz0CtrlAxiBReady;
sGtwiz0CtrlAxiARAddr <= sGtwiz0CtrlAxiARAddr;
sGtwiz0CtrlAxiARValid <= sGtwiz0CtrlAxiARValid;
sGtwiz0CtrlAxiARReady <= sGtwiz0CtrlAxiARReady;
sGtwiz0CtrlAxiRData <= sGtwiz0CtrlAxiRData;
sGtwiz0CtrlAxiRResp <= sGtwiz0CtrlAxiRResp;
sGtwiz0CtrlAxiRValid <= sGtwiz0CtrlAxiRValid;
sGtwiz0CtrlAxiRReady <= sGtwiz0CtrlAxiRReady;
sGtwiz0DrpChAxiAWAddr <= sGtwiz0DrpChAxiAWAddr;
sGtwiz0DrpChAxiAWValid <= sGtwiz0DrpChAxiAWValid;
sGtwiz0DrpChAxiAWReady <= sGtwiz0DrpChAxiAWReady;
sGtwiz0DrpChAxiWData <= sGtwiz0DrpChAxiWData;
sGtwiz0DrpChAxiWStrb <= sGtwiz0DrpChAxiWStrb;
sGtwiz0DrpChAxiWValid <= sGtwiz0DrpChAxiWValid;
sGtwiz0DrpChAxiWReady <= sGtwiz0DrpChAxiWReady;
sGtwiz0DrpChAxiBResp <= sGtwiz0DrpChAxiBResp;
sGtwiz0DrpChAxiBValid <= sGtwiz0DrpChAxiBValid;
sGtwiz0DrpChAxiBReady <= sGtwiz0DrpChAxiBReady;
sGtwiz0DrpChAxiARAddr <= sGtwiz0DrpChAxiARAddr;
sGtwiz0DrpChAxiARValid <= sGtwiz0DrpChAxiARValid;
sGtwiz0DrpChAxiARReady <= sGtwiz0DrpChAxiARReady;
sGtwiz0DrpChAxiRData <= sGtwiz0DrpChAxiRData;
sGtwiz0DrpChAxiRResp <= sGtwiz0DrpChAxiRResp;
sGtwiz0DrpChAxiRValid <= sGtwiz0DrpChAxiRValid;
sGtwiz0DrpChAxiRReady <= sGtwiz0DrpChAxiRReady;
UserClkPort1 <= UserClkPort1;
aPort1PmaInit <= aPort1PmaInit;
aPort1ResetPb <= aPort1ResetPb;
uPort1AxiTxTData0 <= uPort1AxiTxTData0;
uPort1AxiTxTData1 <= uPort1AxiTxTData1;
uPort1AxiTxTData2 <= uPort1AxiTxTData2;
uPort1AxiTxTData3 <= uPort1AxiTxTData3;
uPort1AxiTxTKeep <= uPort1AxiTxTKeep;
uPort1AxiTxTLast <= uPort1AxiTxTLast;
uPort1AxiTxTValid <= uPort1AxiTxTValid;
uPort1AxiTxTReady <= uPort1AxiTxTReady;
uPort1AxiRxTData0 <= uPort1AxiRxTData0;
uPort1AxiRxTData1 <= uPort1AxiRxTData1;
uPort1AxiRxTData2 <= uPort1AxiRxTData2;
uPort1AxiRxTData3 <= uPort1AxiRxTData3;
uPort1AxiRxTKeep <= uPort1AxiRxTKeep;
uPort1AxiRxTLast <= uPort1AxiRxTLast;
uPort1AxiRxTValid <= uPort1AxiRxTValid;
uPort1AxiNfcTValid <= uPort1AxiNfcTValid;
uPort1AxiNfcTData <= uPort1AxiNfcTData;
uPort1AxiNfcTReady <= uPort1AxiNfcTReady;
uPort1HardError <= uPort1HardError;
uPort1SoftError <= uPort1SoftError;
uPort1LaneUp <= uPort1LaneUp;
uPort1ChannelUp <= uPort1ChannelUp;
uPort1SysResetOut <= uPort1SysResetOut;
uPort1MmcmNotLockOut <= uPort1MmcmNotLockOut;
uPort1CrcPassFail_n <= uPort1CrcPassFail_n;
uPort1CrcValid <= uPort1CrcValid;
iPort1LinkResetOut <= iPort1LinkResetOut;
sGtwiz1CtrlAxiAWAddr <= sGtwiz1CtrlAxiAWAddr;
sGtwiz1CtrlAxiAWValid <= sGtwiz1CtrlAxiAWValid;
sGtwiz1CtrlAxiAWReady <= sGtwiz1CtrlAxiAWReady;
sGtwiz1CtrlAxiWData <= sGtwiz1CtrlAxiWData;
sGtwiz1CtrlAxiWStrb <= sGtwiz1CtrlAxiWStrb;
sGtwiz1CtrlAxiWValid <= sGtwiz1CtrlAxiWValid;
sGtwiz1CtrlAxiWReady <= sGtwiz1CtrlAxiWReady;
sGtwiz1CtrlAxiBResp <= sGtwiz1CtrlAxiBResp;
sGtwiz1CtrlAxiBValid <= sGtwiz1CtrlAxiBValid;
sGtwiz1CtrlAxiBReady <= sGtwiz1CtrlAxiBReady;
sGtwiz1CtrlAxiARAddr <= sGtwiz1CtrlAxiARAddr;
sGtwiz1CtrlAxiARValid <= sGtwiz1CtrlAxiARValid;
sGtwiz1CtrlAxiARReady <= sGtwiz1CtrlAxiARReady;
sGtwiz1CtrlAxiRData <= sGtwiz1CtrlAxiRData;
sGtwiz1CtrlAxiRResp <= sGtwiz1CtrlAxiRResp;
sGtwiz1CtrlAxiRValid <= sGtwiz1CtrlAxiRValid;
sGtwiz1CtrlAxiRReady <= sGtwiz1CtrlAxiRReady;
sGtwiz1DrpChAxiAWAddr <= sGtwiz1DrpChAxiAWAddr;
sGtwiz1DrpChAxiAWValid <= sGtwiz1DrpChAxiAWValid;
sGtwiz1DrpChAxiAWReady <= sGtwiz1DrpChAxiAWReady;
sGtwiz1DrpChAxiWData <= sGtwiz1DrpChAxiWData;
sGtwiz1DrpChAxiWStrb <= sGtwiz1DrpChAxiWStrb;
sGtwiz1DrpChAxiWValid <= sGtwiz1DrpChAxiWValid;
sGtwiz1DrpChAxiWReady <= sGtwiz1DrpChAxiWReady;
sGtwiz1DrpChAxiBResp <= sGtwiz1DrpChAxiBResp;
sGtwiz1DrpChAxiBValid <= sGtwiz1DrpChAxiBValid;
sGtwiz1DrpChAxiBReady <= sGtwiz1DrpChAxiBReady;
sGtwiz1DrpChAxiARAddr <= sGtwiz1DrpChAxiARAddr;
sGtwiz1DrpChAxiARValid <= sGtwiz1DrpChAxiARValid;
sGtwiz1DrpChAxiARReady <= sGtwiz1DrpChAxiARReady;
sGtwiz1DrpChAxiRData <= sGtwiz1DrpChAxiRData;
sGtwiz1DrpChAxiRResp <= sGtwiz1DrpChAxiRResp;
sGtwiz1DrpChAxiRValid <= sGtwiz1DrpChAxiRValid;
sGtwiz1DrpChAxiRReady <= sGtwiz1DrpChAxiRReady;
UserClkPort2 <= UserClkPort2;
aPort2PmaInit <= aPort2PmaInit;
aPort2ResetPb <= aPort2ResetPb;
uPort2AxiTxTData0 <= uPort2AxiTxTData0;
uPort2AxiTxTData1 <= uPort2AxiTxTData1;
uPort2AxiTxTData2 <= uPort2AxiTxTData2;
uPort2AxiTxTData3 <= uPort2AxiTxTData3;
uPort2AxiTxTKeep <= uPort2AxiTxTKeep;
uPort2AxiTxTLast <= uPort2AxiTxTLast;
uPort2AxiTxTValid <= uPort2AxiTxTValid;
uPort2AxiTxTReady <= uPort2AxiTxTReady;
uPort2AxiRxTData0 <= uPort2AxiRxTData0;
uPort2AxiRxTData1 <= uPort2AxiRxTData1;
uPort2AxiRxTData2 <= uPort2AxiRxTData2;
uPort2AxiRxTData3 <= uPort2AxiRxTData3;
uPort2AxiRxTKeep <= uPort2AxiRxTKeep;
uPort2AxiRxTLast <= uPort2AxiRxTLast;
uPort2AxiRxTValid <= uPort2AxiRxTValid;
uPort2AxiNfcTValid <= uPort2AxiNfcTValid;
uPort2AxiNfcTData <= uPort2AxiNfcTData;
uPort2AxiNfcTReady <= uPort2AxiNfcTReady;
uPort2HardError <= uPort2HardError;
uPort2SoftError <= uPort2SoftError;
uPort2LaneUp <= uPort2LaneUp;
uPort2ChannelUp <= uPort2ChannelUp;
uPort2SysResetOut <= uPort2SysResetOut;
uPort2MmcmNotLockOut <= uPort2MmcmNotLockOut;
uPort2CrcPassFail_n <= uPort2CrcPassFail_n;
uPort2CrcValid <= uPort2CrcValid;
iPort2LinkResetOut <= iPort2LinkResetOut;
sGtwiz2CtrlAxiAWAddr <= sGtwiz2CtrlAxiAWAddr;
sGtwiz2CtrlAxiAWValid <= sGtwiz2CtrlAxiAWValid;
sGtwiz2CtrlAxiAWReady <= sGtwiz2CtrlAxiAWReady;
sGtwiz2CtrlAxiWData <= sGtwiz2CtrlAxiWData;
sGtwiz2CtrlAxiWStrb <= sGtwiz2CtrlAxiWStrb;
sGtwiz2CtrlAxiWValid <= sGtwiz2CtrlAxiWValid;
sGtwiz2CtrlAxiWReady <= sGtwiz2CtrlAxiWReady;
sGtwiz2CtrlAxiBResp <= sGtwiz2CtrlAxiBResp;
sGtwiz2CtrlAxiBValid <= sGtwiz2CtrlAxiBValid;
sGtwiz2CtrlAxiBReady <= sGtwiz2CtrlAxiBReady;
sGtwiz2CtrlAxiARAddr <= sGtwiz2CtrlAxiARAddr;
sGtwiz2CtrlAxiARValid <= sGtwiz2CtrlAxiARValid;
sGtwiz2CtrlAxiARReady <= sGtwiz2CtrlAxiARReady;
sGtwiz2CtrlAxiRData <= sGtwiz2CtrlAxiRData;
sGtwiz2CtrlAxiRResp <= sGtwiz2CtrlAxiRResp;
sGtwiz2CtrlAxiRValid <= sGtwiz2CtrlAxiRValid;
sGtwiz2CtrlAxiRReady <= sGtwiz2CtrlAxiRReady;
sGtwiz2DrpChAxiAWAddr <= sGtwiz2DrpChAxiAWAddr;
sGtwiz2DrpChAxiAWValid <= sGtwiz2DrpChAxiAWValid;
sGtwiz2DrpChAxiAWReady <= sGtwiz2DrpChAxiAWReady;
sGtwiz2DrpChAxiWData <= sGtwiz2DrpChAxiWData;
sGtwiz2DrpChAxiWStrb <= sGtwiz2DrpChAxiWStrb;
sGtwiz2DrpChAxiWValid <= sGtwiz2DrpChAxiWValid;
sGtwiz2DrpChAxiWReady <= sGtwiz2DrpChAxiWReady;
sGtwiz2DrpChAxiBResp <= sGtwiz2DrpChAxiBResp;
sGtwiz2DrpChAxiBValid <= sGtwiz2DrpChAxiBValid;
sGtwiz2DrpChAxiBReady <= sGtwiz2DrpChAxiBReady;
sGtwiz2DrpChAxiARAddr <= sGtwiz2DrpChAxiARAddr;
sGtwiz2DrpChAxiARValid <= sGtwiz2DrpChAxiARValid;
sGtwiz2DrpChAxiARReady <= sGtwiz2DrpChAxiARReady;
sGtwiz2DrpChAxiRData <= sGtwiz2DrpChAxiRData;
sGtwiz2DrpChAxiRResp <= sGtwiz2DrpChAxiRResp;
sGtwiz2DrpChAxiRValid <= sGtwiz2DrpChAxiRValid;
sGtwiz2DrpChAxiRReady <= sGtwiz2DrpChAxiRReady;
UserClkPort3 <= UserClkPort3;
aPort3PmaInit <= aPort3PmaInit;
aPort3ResetPb <= aPort3ResetPb;
uPort3AxiTxTData0 <= uPort3AxiTxTData0;
uPort3AxiTxTData1 <= uPort3AxiTxTData1;
uPort3AxiTxTData2 <= uPort3AxiTxTData2;
uPort3AxiTxTData3 <= uPort3AxiTxTData3;
uPort3AxiTxTKeep <= uPort3AxiTxTKeep;
uPort3AxiTxTLast <= uPort3AxiTxTLast;
uPort3AxiTxTValid <= uPort3AxiTxTValid;
uPort3AxiTxTReady <= uPort3AxiTxTReady;
uPort3AxiRxTData0 <= uPort3AxiRxTData0;
uPort3AxiRxTData1 <= uPort3AxiRxTData1;
uPort3AxiRxTData2 <= uPort3AxiRxTData2;
uPort3AxiRxTData3 <= uPort3AxiRxTData3;
uPort3AxiRxTKeep <= uPort3AxiRxTKeep;
uPort3AxiRxTLast <= uPort3AxiRxTLast;
uPort3AxiRxTValid <= uPort3AxiRxTValid;
uPort3AxiNfcTValid <= uPort3AxiNfcTValid;
uPort3AxiNfcTData <= uPort3AxiNfcTData;
uPort3AxiNfcTReady <= uPort3AxiNfcTReady;
uPort3HardError <= uPort3HardError;
uPort3SoftError <= uPort3SoftError;
uPort3LaneUp <= uPort3LaneUp;
uPort3ChannelUp <= uPort3ChannelUp;
uPort3SysResetOut <= uPort3SysResetOut;
uPort3MmcmNotLockOut <= uPort3MmcmNotLockOut;
uPort3CrcPassFail_n <= uPort3CrcPassFail_n;
uPort3CrcValid <= uPort3CrcValid;
iPort3LinkResetOut <= iPort3LinkResetOut;
sGtwiz3CtrlAxiAWAddr <= sGtwiz3CtrlAxiAWAddr;
sGtwiz3CtrlAxiAWValid <= sGtwiz3CtrlAxiAWValid;
sGtwiz3CtrlAxiAWReady <= sGtwiz3CtrlAxiAWReady;
sGtwiz3CtrlAxiWData <= sGtwiz3CtrlAxiWData;
sGtwiz3CtrlAxiWStrb <= sGtwiz3CtrlAxiWStrb;
sGtwiz3CtrlAxiWValid <= sGtwiz3CtrlAxiWValid;
sGtwiz3CtrlAxiWReady <= sGtwiz3CtrlAxiWReady;
sGtwiz3CtrlAxiBResp <= sGtwiz3CtrlAxiBResp;
sGtwiz3CtrlAxiBValid <= sGtwiz3CtrlAxiBValid;
sGtwiz3CtrlAxiBReady <= sGtwiz3CtrlAxiBReady;
sGtwiz3CtrlAxiARAddr <= sGtwiz3CtrlAxiARAddr;
sGtwiz3CtrlAxiARValid <= sGtwiz3CtrlAxiARValid;
sGtwiz3CtrlAxiARReady <= sGtwiz3CtrlAxiARReady;
sGtwiz3CtrlAxiRData <= sGtwiz3CtrlAxiRData;
sGtwiz3CtrlAxiRResp <= sGtwiz3CtrlAxiRResp;
sGtwiz3CtrlAxiRValid <= sGtwiz3CtrlAxiRValid;
sGtwiz3CtrlAxiRReady <= sGtwiz3CtrlAxiRReady;
sGtwiz3DrpChAxiAWAddr <= sGtwiz3DrpChAxiAWAddr;
sGtwiz3DrpChAxiAWValid <= sGtwiz3DrpChAxiAWValid;
sGtwiz3DrpChAxiAWReady <= sGtwiz3DrpChAxiAWReady;
sGtwiz3DrpChAxiWData <= sGtwiz3DrpChAxiWData;
sGtwiz3DrpChAxiWStrb <= sGtwiz3DrpChAxiWStrb;
sGtwiz3DrpChAxiWValid <= sGtwiz3DrpChAxiWValid;
sGtwiz3DrpChAxiWReady <= sGtwiz3DrpChAxiWReady;
sGtwiz3DrpChAxiBResp <= sGtwiz3DrpChAxiBResp;
sGtwiz3DrpChAxiBValid <= sGtwiz3DrpChAxiBValid;
sGtwiz3DrpChAxiBReady <= sGtwiz3DrpChAxiBReady;
sGtwiz3DrpChAxiARAddr <= sGtwiz3DrpChAxiARAddr;
sGtwiz3DrpChAxiARValid <= sGtwiz3DrpChAxiARValid;
sGtwiz3DrpChAxiARReady <= sGtwiz3DrpChAxiARReady;
sGtwiz3DrpChAxiRData <= sGtwiz3DrpChAxiRData;
sGtwiz3DrpChAxiRResp <= sGtwiz3DrpChAxiRResp;
sGtwiz3DrpChAxiRValid <= sGtwiz3DrpChAxiRValid;
sGtwiz3DrpChAxiRReady <= sGtwiz3DrpChAxiRReady;
UserClkPort4 <= UserClkPort4;
aPort4PmaInit <= aPort4PmaInit;
aPort4ResetPb <= aPort4ResetPb;
uPort4AxiTxTData0 <= uPort4AxiTxTData0;
uPort4AxiTxTData1 <= uPort4AxiTxTData1;
uPort4AxiTxTData2 <= uPort4AxiTxTData2;
uPort4AxiTxTData3 <= uPort4AxiTxTData3;
uPort4AxiTxTKeep <= uPort4AxiTxTKeep;
uPort4AxiTxTLast <= uPort4AxiTxTLast;
uPort4AxiTxTValid <= uPort4AxiTxTValid;
uPort4AxiTxTReady <= uPort4AxiTxTReady;
uPort4AxiRxTData0 <= uPort4AxiRxTData0;
uPort4AxiRxTData1 <= uPort4AxiRxTData1;
uPort4AxiRxTData2 <= uPort4AxiRxTData2;
uPort4AxiRxTData3 <= uPort4AxiRxTData3;
uPort4AxiRxTKeep <= uPort4AxiRxTKeep;
uPort4AxiRxTLast <= uPort4AxiRxTLast;
uPort4AxiRxTValid <= uPort4AxiRxTValid;
uPort4AxiNfcTValid <= uPort4AxiNfcTValid;
uPort4AxiNfcTData <= uPort4AxiNfcTData;
uPort4AxiNfcTReady <= uPort4AxiNfcTReady;
uPort4HardError <= uPort4HardError;
uPort4SoftError <= uPort4SoftError;
uPort4LaneUp <= uPort4LaneUp;
uPort4ChannelUp <= uPort4ChannelUp;
uPort4SysResetOut <= uPort4SysResetOut;
uPort4MmcmNotLockOut <= uPort4MmcmNotLockOut;
uPort4CrcPassFail_n <= uPort4CrcPassFail_n;
uPort4CrcValid <= uPort4CrcValid;
iPort4LinkResetOut <= iPort4LinkResetOut;
sGtwiz4CtrlAxiAWAddr <= sGtwiz4CtrlAxiAWAddr;
sGtwiz4CtrlAxiAWValid <= sGtwiz4CtrlAxiAWValid;
sGtwiz4CtrlAxiAWReady <= sGtwiz4CtrlAxiAWReady;
sGtwiz4CtrlAxiWData <= sGtwiz4CtrlAxiWData;
sGtwiz4CtrlAxiWStrb <= sGtwiz4CtrlAxiWStrb;
sGtwiz4CtrlAxiWValid <= sGtwiz4CtrlAxiWValid;
sGtwiz4CtrlAxiWReady <= sGtwiz4CtrlAxiWReady;
sGtwiz4CtrlAxiBResp <= sGtwiz4CtrlAxiBResp;
sGtwiz4CtrlAxiBValid <= sGtwiz4CtrlAxiBValid;
sGtwiz4CtrlAxiBReady <= sGtwiz4CtrlAxiBReady;
sGtwiz4CtrlAxiARAddr <= sGtwiz4CtrlAxiARAddr;
sGtwiz4CtrlAxiARValid <= sGtwiz4CtrlAxiARValid;
sGtwiz4CtrlAxiARReady <= sGtwiz4CtrlAxiARReady;
sGtwiz4CtrlAxiRData <= sGtwiz4CtrlAxiRData;
sGtwiz4CtrlAxiRResp <= sGtwiz4CtrlAxiRResp;
sGtwiz4CtrlAxiRValid <= sGtwiz4CtrlAxiRValid;
sGtwiz4CtrlAxiRReady <= sGtwiz4CtrlAxiRReady;
sGtwiz4DrpChAxiAWAddr <= sGtwiz4DrpChAxiAWAddr;
sGtwiz4DrpChAxiAWValid <= sGtwiz4DrpChAxiAWValid;
sGtwiz4DrpChAxiAWReady <= sGtwiz4DrpChAxiAWReady;
sGtwiz4DrpChAxiWData <= sGtwiz4DrpChAxiWData;
sGtwiz4DrpChAxiWStrb <= sGtwiz4DrpChAxiWStrb;
sGtwiz4DrpChAxiWValid <= sGtwiz4DrpChAxiWValid;
sGtwiz4DrpChAxiWReady <= sGtwiz4DrpChAxiWReady;
sGtwiz4DrpChAxiBResp <= sGtwiz4DrpChAxiBResp;
sGtwiz4DrpChAxiBValid <= sGtwiz4DrpChAxiBValid;
sGtwiz4DrpChAxiBReady <= sGtwiz4DrpChAxiBReady;
sGtwiz4DrpChAxiARAddr <= sGtwiz4DrpChAxiARAddr;
sGtwiz4DrpChAxiARValid <= sGtwiz4DrpChAxiARValid;
sGtwiz4DrpChAxiARReady <= sGtwiz4DrpChAxiARReady;
sGtwiz4DrpChAxiRData <= sGtwiz4DrpChAxiRData;
sGtwiz4DrpChAxiRResp <= sGtwiz4DrpChAxiRResp;
sGtwiz4DrpChAxiRValid <= sGtwiz4DrpChAxiRValid;
sGtwiz4DrpChAxiRReady <= sGtwiz4DrpChAxiRReady;
UserClkPort5 <= UserClkPort5;
aPort5PmaInit <= aPort5PmaInit;
aPort5ResetPb <= aPort5ResetPb;
uPort5AxiTxTData0 <= uPort5AxiTxTData0;
uPort5AxiTxTData1 <= uPort5AxiTxTData1;
uPort5AxiTxTData2 <= uPort5AxiTxTData2;
uPort5AxiTxTData3 <= uPort5AxiTxTData3;
uPort5AxiTxTKeep <= uPort5AxiTxTKeep;
uPort5AxiTxTLast <= uPort5AxiTxTLast;
uPort5AxiTxTValid <= uPort5AxiTxTValid;
uPort5AxiTxTReady <= uPort5AxiTxTReady;
uPort5AxiRxTData0 <= uPort5AxiRxTData0;
uPort5AxiRxTData1 <= uPort5AxiRxTData1;
uPort5AxiRxTData2 <= uPort5AxiRxTData2;
uPort5AxiRxTData3 <= uPort5AxiRxTData3;
uPort5AxiRxTKeep <= uPort5AxiRxTKeep;
uPort5AxiRxTLast <= uPort5AxiRxTLast;
uPort5AxiRxTValid <= uPort5AxiRxTValid;
uPort5AxiNfcTValid <= uPort5AxiNfcTValid;
uPort5AxiNfcTData <= uPort5AxiNfcTData;
uPort5AxiNfcTReady <= uPort5AxiNfcTReady;
uPort5HardError <= uPort5HardError;
uPort5SoftError <= uPort5SoftError;
uPort5LaneUp <= uPort5LaneUp;
uPort5ChannelUp <= uPort5ChannelUp;
uPort5SysResetOut <= uPort5SysResetOut;
uPort5MmcmNotLockOut <= uPort5MmcmNotLockOut;
uPort5CrcPassFail_n <= uPort5CrcPassFail_n;
uPort5CrcValid <= uPort5CrcValid;
iPort5LinkResetOut <= iPort5LinkResetOut;
sGtwiz5CtrlAxiAWAddr <= sGtwiz5CtrlAxiAWAddr;
sGtwiz5CtrlAxiAWValid <= sGtwiz5CtrlAxiAWValid;
sGtwiz5CtrlAxiAWReady <= sGtwiz5CtrlAxiAWReady;
sGtwiz5CtrlAxiWData <= sGtwiz5CtrlAxiWData;
sGtwiz5CtrlAxiWStrb <= sGtwiz5CtrlAxiWStrb;
sGtwiz5CtrlAxiWValid <= sGtwiz5CtrlAxiWValid;
sGtwiz5CtrlAxiWReady <= sGtwiz5CtrlAxiWReady;
sGtwiz5CtrlAxiBResp <= sGtwiz5CtrlAxiBResp;
sGtwiz5CtrlAxiBValid <= sGtwiz5CtrlAxiBValid;
sGtwiz5CtrlAxiBReady <= sGtwiz5CtrlAxiBReady;
sGtwiz5CtrlAxiARAddr <= sGtwiz5CtrlAxiARAddr;
sGtwiz5CtrlAxiARValid <= sGtwiz5CtrlAxiARValid;
sGtwiz5CtrlAxiARReady <= sGtwiz5CtrlAxiARReady;
sGtwiz5CtrlAxiRData <= sGtwiz5CtrlAxiRData;
sGtwiz5CtrlAxiRResp <= sGtwiz5CtrlAxiRResp;
sGtwiz5CtrlAxiRValid <= sGtwiz5CtrlAxiRValid;
sGtwiz5CtrlAxiRReady <= sGtwiz5CtrlAxiRReady;
sGtwiz5DrpChAxiAWAddr <= sGtwiz5DrpChAxiAWAddr;
sGtwiz5DrpChAxiAWValid <= sGtwiz5DrpChAxiAWValid;
sGtwiz5DrpChAxiAWReady <= sGtwiz5DrpChAxiAWReady;
sGtwiz5DrpChAxiWData <= sGtwiz5DrpChAxiWData;
sGtwiz5DrpChAxiWStrb <= sGtwiz5DrpChAxiWStrb;
sGtwiz5DrpChAxiWValid <= sGtwiz5DrpChAxiWValid;
sGtwiz5DrpChAxiWReady <= sGtwiz5DrpChAxiWReady;
sGtwiz5DrpChAxiBResp <= sGtwiz5DrpChAxiBResp;
sGtwiz5DrpChAxiBValid <= sGtwiz5DrpChAxiBValid;
sGtwiz5DrpChAxiBReady <= sGtwiz5DrpChAxiBReady;
sGtwiz5DrpChAxiARAddr <= sGtwiz5DrpChAxiARAddr;
sGtwiz5DrpChAxiARValid <= sGtwiz5DrpChAxiARValid;
sGtwiz5DrpChAxiARReady <= sGtwiz5DrpChAxiARReady;
sGtwiz5DrpChAxiRData <= sGtwiz5DrpChAxiRData;
sGtwiz5DrpChAxiRResp <= sGtwiz5DrpChAxiRResp;
sGtwiz5DrpChAxiRValid <= sGtwiz5DrpChAxiRValid;
sGtwiz5DrpChAxiRReady <= sGtwiz5DrpChAxiRReady;
UserClkPort6 <= UserClkPort6;
aPort6PmaInit <= aPort6PmaInit;
aPort6ResetPb <= aPort6ResetPb;
uPort6AxiTxTData0 <= uPort6AxiTxTData0;
uPort6AxiTxTData1 <= uPort6AxiTxTData1;
uPort6AxiTxTData2 <= uPort6AxiTxTData2;
uPort6AxiTxTData3 <= uPort6AxiTxTData3;
uPort6AxiTxTKeep <= uPort6AxiTxTKeep;
uPort6AxiTxTLast <= uPort6AxiTxTLast;
uPort6AxiTxTValid <= uPort6AxiTxTValid;
uPort6AxiTxTReady <= uPort6AxiTxTReady;
uPort6AxiRxTData0 <= uPort6AxiRxTData0;
uPort6AxiRxTData1 <= uPort6AxiRxTData1;
uPort6AxiRxTData2 <= uPort6AxiRxTData2;
uPort6AxiRxTData3 <= uPort6AxiRxTData3;
uPort6AxiRxTKeep <= uPort6AxiRxTKeep;
uPort6AxiRxTLast <= uPort6AxiRxTLast;
uPort6AxiRxTValid <= uPort6AxiRxTValid;
uPort6AxiNfcTValid <= uPort6AxiNfcTValid;
uPort6AxiNfcTData <= uPort6AxiNfcTData;
uPort6AxiNfcTReady <= uPort6AxiNfcTReady;
uPort6HardError <= uPort6HardError;
uPort6SoftError <= uPort6SoftError;
uPort6LaneUp <= uPort6LaneUp;
uPort6ChannelUp <= uPort6ChannelUp;
uPort6SysResetOut <= uPort6SysResetOut;
uPort6MmcmNotLockOut <= uPort6MmcmNotLockOut;
uPort6CrcPassFail_n <= uPort6CrcPassFail_n;
uPort6CrcValid <= uPort6CrcValid;
iPort6LinkResetOut <= iPort6LinkResetOut;
sGtwiz6CtrlAxiAWAddr <= sGtwiz6CtrlAxiAWAddr;
sGtwiz6CtrlAxiAWValid <= sGtwiz6CtrlAxiAWValid;
sGtwiz6CtrlAxiAWReady <= sGtwiz6CtrlAxiAWReady;
sGtwiz6CtrlAxiWData <= sGtwiz6CtrlAxiWData;
sGtwiz6CtrlAxiWStrb <= sGtwiz6CtrlAxiWStrb;
sGtwiz6CtrlAxiWValid <= sGtwiz6CtrlAxiWValid;
sGtwiz6CtrlAxiWReady <= sGtwiz6CtrlAxiWReady;
sGtwiz6CtrlAxiBResp <= sGtwiz6CtrlAxiBResp;
sGtwiz6CtrlAxiBValid <= sGtwiz6CtrlAxiBValid;
sGtwiz6CtrlAxiBReady <= sGtwiz6CtrlAxiBReady;
sGtwiz6CtrlAxiARAddr <= sGtwiz6CtrlAxiARAddr;
sGtwiz6CtrlAxiARValid <= sGtwiz6CtrlAxiARValid;
sGtwiz6CtrlAxiARReady <= sGtwiz6CtrlAxiARReady;
sGtwiz6CtrlAxiRData <= sGtwiz6CtrlAxiRData;
sGtwiz6CtrlAxiRResp <= sGtwiz6CtrlAxiRResp;
sGtwiz6CtrlAxiRValid <= sGtwiz6CtrlAxiRValid;
sGtwiz6CtrlAxiRReady <= sGtwiz6CtrlAxiRReady;
sGtwiz6DrpChAxiAWAddr <= sGtwiz6DrpChAxiAWAddr;
sGtwiz6DrpChAxiAWValid <= sGtwiz6DrpChAxiAWValid;
sGtwiz6DrpChAxiAWReady <= sGtwiz6DrpChAxiAWReady;
sGtwiz6DrpChAxiWData <= sGtwiz6DrpChAxiWData;
sGtwiz6DrpChAxiWStrb <= sGtwiz6DrpChAxiWStrb;
sGtwiz6DrpChAxiWValid <= sGtwiz6DrpChAxiWValid;
sGtwiz6DrpChAxiWReady <= sGtwiz6DrpChAxiWReady;
sGtwiz6DrpChAxiBResp <= sGtwiz6DrpChAxiBResp;
sGtwiz6DrpChAxiBValid <= sGtwiz6DrpChAxiBValid;
sGtwiz6DrpChAxiBReady <= sGtwiz6DrpChAxiBReady;
sGtwiz6DrpChAxiARAddr <= sGtwiz6DrpChAxiARAddr;
sGtwiz6DrpChAxiARValid <= sGtwiz6DrpChAxiARValid;
sGtwiz6DrpChAxiARReady <= sGtwiz6DrpChAxiARReady;
sGtwiz6DrpChAxiRData <= sGtwiz6DrpChAxiRData;
sGtwiz6DrpChAxiRResp <= sGtwiz6DrpChAxiRResp;
sGtwiz6DrpChAxiRValid <= sGtwiz6DrpChAxiRValid;
sGtwiz6DrpChAxiRReady <= sGtwiz6DrpChAxiRReady;
UserClkPort7 <= UserClkPort7;
aPort7PmaInit <= aPort7PmaInit;
aPort7ResetPb <= aPort7ResetPb;
uPort7AxiTxTData0 <= uPort7AxiTxTData0;
uPort7AxiTxTData1 <= uPort7AxiTxTData1;
uPort7AxiTxTData2 <= uPort7AxiTxTData2;
uPort7AxiTxTData3 <= uPort7AxiTxTData3;
uPort7AxiTxTKeep <= uPort7AxiTxTKeep;
uPort7AxiTxTLast <= uPort7AxiTxTLast;
uPort7AxiTxTValid <= uPort7AxiTxTValid;
uPort7AxiTxTReady <= uPort7AxiTxTReady;
uPort7AxiRxTData0 <= uPort7AxiRxTData0;
uPort7AxiRxTData1 <= uPort7AxiRxTData1;
uPort7AxiRxTData2 <= uPort7AxiRxTData2;
uPort7AxiRxTData3 <= uPort7AxiRxTData3;
uPort7AxiRxTKeep <= uPort7AxiRxTKeep;
uPort7AxiRxTLast <= uPort7AxiRxTLast;
uPort7AxiRxTValid <= uPort7AxiRxTValid;
uPort7AxiNfcTValid <= uPort7AxiNfcTValid;
uPort7AxiNfcTData <= uPort7AxiNfcTData;
uPort7AxiNfcTReady <= uPort7AxiNfcTReady;
uPort7HardError <= uPort7HardError;
uPort7SoftError <= uPort7SoftError;
uPort7LaneUp <= uPort7LaneUp;
uPort7ChannelUp <= uPort7ChannelUp;
uPort7SysResetOut <= uPort7SysResetOut;
uPort7MmcmNotLockOut <= uPort7MmcmNotLockOut;
uPort7CrcPassFail_n <= uPort7CrcPassFail_n;
uPort7CrcValid <= uPort7CrcValid;
iPort7LinkResetOut <= iPort7LinkResetOut;
sGtwiz7CtrlAxiAWAddr <= sGtwiz7CtrlAxiAWAddr;
sGtwiz7CtrlAxiAWValid <= sGtwiz7CtrlAxiAWValid;
sGtwiz7CtrlAxiAWReady <= sGtwiz7CtrlAxiAWReady;
sGtwiz7CtrlAxiWData <= sGtwiz7CtrlAxiWData;
sGtwiz7CtrlAxiWStrb <= sGtwiz7CtrlAxiWStrb;
sGtwiz7CtrlAxiWValid <= sGtwiz7CtrlAxiWValid;
sGtwiz7CtrlAxiWReady <= sGtwiz7CtrlAxiWReady;
sGtwiz7CtrlAxiBResp <= sGtwiz7CtrlAxiBResp;
sGtwiz7CtrlAxiBValid <= sGtwiz7CtrlAxiBValid;
sGtwiz7CtrlAxiBReady <= sGtwiz7CtrlAxiBReady;
sGtwiz7CtrlAxiARAddr <= sGtwiz7CtrlAxiARAddr;
sGtwiz7CtrlAxiARValid <= sGtwiz7CtrlAxiARValid;
sGtwiz7CtrlAxiARReady <= sGtwiz7CtrlAxiARReady;
sGtwiz7CtrlAxiRData <= sGtwiz7CtrlAxiRData;
sGtwiz7CtrlAxiRResp <= sGtwiz7CtrlAxiRResp;
sGtwiz7CtrlAxiRValid <= sGtwiz7CtrlAxiRValid;
sGtwiz7CtrlAxiRReady <= sGtwiz7CtrlAxiRReady;
sGtwiz7DrpChAxiAWAddr <= sGtwiz7DrpChAxiAWAddr;
sGtwiz7DrpChAxiAWValid <= sGtwiz7DrpChAxiAWValid;
sGtwiz7DrpChAxiAWReady <= sGtwiz7DrpChAxiAWReady;
sGtwiz7DrpChAxiWData <= sGtwiz7DrpChAxiWData;
sGtwiz7DrpChAxiWStrb <= sGtwiz7DrpChAxiWStrb;
sGtwiz7DrpChAxiWValid <= sGtwiz7DrpChAxiWValid;
sGtwiz7DrpChAxiWReady <= sGtwiz7DrpChAxiWReady;
sGtwiz7DrpChAxiBResp <= sGtwiz7DrpChAxiBResp;
sGtwiz7DrpChAxiBValid <= sGtwiz7DrpChAxiBValid;
sGtwiz7DrpChAxiBReady <= sGtwiz7DrpChAxiBReady;
sGtwiz7DrpChAxiARAddr <= sGtwiz7DrpChAxiARAddr;
sGtwiz7DrpChAxiARValid <= sGtwiz7DrpChAxiARValid;
sGtwiz7DrpChAxiARReady <= sGtwiz7DrpChAxiARReady;
sGtwiz7DrpChAxiRData <= sGtwiz7DrpChAxiRData;
sGtwiz7DrpChAxiRResp <= sGtwiz7DrpChAxiRResp;
sGtwiz7DrpChAxiRValid <= sGtwiz7DrpChAxiRValid;
sGtwiz7DrpChAxiRReady <= sGtwiz7DrpChAxiRReady;
UserClkPort8 <= UserClkPort8;
aPort8PmaInit <= aPort8PmaInit;
aPort8ResetPb <= aPort8ResetPb;
uPort8AxiTxTData0 <= uPort8AxiTxTData0;
uPort8AxiTxTData1 <= uPort8AxiTxTData1;
uPort8AxiTxTData2 <= uPort8AxiTxTData2;
uPort8AxiTxTData3 <= uPort8AxiTxTData3;
uPort8AxiTxTKeep <= uPort8AxiTxTKeep;
uPort8AxiTxTLast <= uPort8AxiTxTLast;
uPort8AxiTxTValid <= uPort8AxiTxTValid;
uPort8AxiTxTReady <= uPort8AxiTxTReady;
uPort8AxiRxTData0 <= uPort8AxiRxTData0;
uPort8AxiRxTData1 <= uPort8AxiRxTData1;
uPort8AxiRxTData2 <= uPort8AxiRxTData2;
uPort8AxiRxTData3 <= uPort8AxiRxTData3;
uPort8AxiRxTKeep <= uPort8AxiRxTKeep;
uPort8AxiRxTLast <= uPort8AxiRxTLast;
uPort8AxiRxTValid <= uPort8AxiRxTValid;
uPort8AxiNfcTValid <= uPort8AxiNfcTValid;
uPort8AxiNfcTData <= uPort8AxiNfcTData;
uPort8AxiNfcTReady <= uPort8AxiNfcTReady;
uPort8HardError <= uPort8HardError;
uPort8SoftError <= uPort8SoftError;
uPort8LaneUp <= uPort8LaneUp;
uPort8ChannelUp <= uPort8ChannelUp;
uPort8SysResetOut <= uPort8SysResetOut;
uPort8MmcmNotLockOut <= uPort8MmcmNotLockOut;
uPort8CrcPassFail_n <= uPort8CrcPassFail_n;
uPort8CrcValid <= uPort8CrcValid;
iPort8LinkResetOut <= iPort8LinkResetOut;
sGtwiz8CtrlAxiAWAddr <= sGtwiz8CtrlAxiAWAddr;
sGtwiz8CtrlAxiAWValid <= sGtwiz8CtrlAxiAWValid;
sGtwiz8CtrlAxiAWReady <= sGtwiz8CtrlAxiAWReady;
sGtwiz8CtrlAxiWData <= sGtwiz8CtrlAxiWData;
sGtwiz8CtrlAxiWStrb <= sGtwiz8CtrlAxiWStrb;
sGtwiz8CtrlAxiWValid <= sGtwiz8CtrlAxiWValid;
sGtwiz8CtrlAxiWReady <= sGtwiz8CtrlAxiWReady;
sGtwiz8CtrlAxiBResp <= sGtwiz8CtrlAxiBResp;
sGtwiz8CtrlAxiBValid <= sGtwiz8CtrlAxiBValid;
sGtwiz8CtrlAxiBReady <= sGtwiz8CtrlAxiBReady;
sGtwiz8CtrlAxiARAddr <= sGtwiz8CtrlAxiARAddr;
sGtwiz8CtrlAxiARValid <= sGtwiz8CtrlAxiARValid;
sGtwiz8CtrlAxiARReady <= sGtwiz8CtrlAxiARReady;
sGtwiz8CtrlAxiRData <= sGtwiz8CtrlAxiRData;
sGtwiz8CtrlAxiRResp <= sGtwiz8CtrlAxiRResp;
sGtwiz8CtrlAxiRValid <= sGtwiz8CtrlAxiRValid;
sGtwiz8CtrlAxiRReady <= sGtwiz8CtrlAxiRReady;
sGtwiz8DrpChAxiAWAddr <= sGtwiz8DrpChAxiAWAddr;
sGtwiz8DrpChAxiAWValid <= sGtwiz8DrpChAxiAWValid;
sGtwiz8DrpChAxiAWReady <= sGtwiz8DrpChAxiAWReady;
sGtwiz8DrpChAxiWData <= sGtwiz8DrpChAxiWData;
sGtwiz8DrpChAxiWStrb <= sGtwiz8DrpChAxiWStrb;
sGtwiz8DrpChAxiWValid <= sGtwiz8DrpChAxiWValid;
sGtwiz8DrpChAxiWReady <= sGtwiz8DrpChAxiWReady;
sGtwiz8DrpChAxiBResp <= sGtwiz8DrpChAxiBResp;
sGtwiz8DrpChAxiBValid <= sGtwiz8DrpChAxiBValid;
sGtwiz8DrpChAxiBReady <= sGtwiz8DrpChAxiBReady;
sGtwiz8DrpChAxiARAddr <= sGtwiz8DrpChAxiARAddr;
sGtwiz8DrpChAxiARValid <= sGtwiz8DrpChAxiARValid;
sGtwiz8DrpChAxiARReady <= sGtwiz8DrpChAxiARReady;
sGtwiz8DrpChAxiRData <= sGtwiz8DrpChAxiRData;
sGtwiz8DrpChAxiRResp <= sGtwiz8DrpChAxiRResp;
sGtwiz8DrpChAxiRValid <= sGtwiz8DrpChAxiRValid;
sGtwiz8DrpChAxiRReady <= sGtwiz8DrpChAxiRReady;
UserClkPort9 <= UserClkPort9;
aPort9PmaInit <= aPort9PmaInit;
aPort9ResetPb <= aPort9ResetPb;
uPort9AxiTxTData0 <= uPort9AxiTxTData0;
uPort9AxiTxTData1 <= uPort9AxiTxTData1;
uPort9AxiTxTData2 <= uPort9AxiTxTData2;
uPort9AxiTxTData3 <= uPort9AxiTxTData3;
uPort9AxiTxTKeep <= uPort9AxiTxTKeep;
uPort9AxiTxTLast <= uPort9AxiTxTLast;
uPort9AxiTxTValid <= uPort9AxiTxTValid;
uPort9AxiTxTReady <= uPort9AxiTxTReady;
uPort9AxiRxTData0 <= uPort9AxiRxTData0;
uPort9AxiRxTData1 <= uPort9AxiRxTData1;
uPort9AxiRxTData2 <= uPort9AxiRxTData2;
uPort9AxiRxTData3 <= uPort9AxiRxTData3;
uPort9AxiRxTKeep <= uPort9AxiRxTKeep;
uPort9AxiRxTLast <= uPort9AxiRxTLast;
uPort9AxiRxTValid <= uPort9AxiRxTValid;
uPort9AxiNfcTValid <= uPort9AxiNfcTValid;
uPort9AxiNfcTData <= uPort9AxiNfcTData;
uPort9AxiNfcTReady <= uPort9AxiNfcTReady;
uPort9HardError <= uPort9HardError;
uPort9SoftError <= uPort9SoftError;
uPort9LaneUp <= uPort9LaneUp;
uPort9ChannelUp <= uPort9ChannelUp;
uPort9SysResetOut <= uPort9SysResetOut;
uPort9MmcmNotLockOut <= uPort9MmcmNotLockOut;
uPort9CrcPassFail_n <= uPort9CrcPassFail_n;
uPort9CrcValid <= uPort9CrcValid;
iPort9LinkResetOut <= iPort9LinkResetOut;
sGtwiz9CtrlAxiAWAddr <= sGtwiz9CtrlAxiAWAddr;
sGtwiz9CtrlAxiAWValid <= sGtwiz9CtrlAxiAWValid;
sGtwiz9CtrlAxiAWReady <= sGtwiz9CtrlAxiAWReady;
sGtwiz9CtrlAxiWData <= sGtwiz9CtrlAxiWData;
sGtwiz9CtrlAxiWStrb <= sGtwiz9CtrlAxiWStrb;
sGtwiz9CtrlAxiWValid <= sGtwiz9CtrlAxiWValid;
sGtwiz9CtrlAxiWReady <= sGtwiz9CtrlAxiWReady;
sGtwiz9CtrlAxiBResp <= sGtwiz9CtrlAxiBResp;
sGtwiz9CtrlAxiBValid <= sGtwiz9CtrlAxiBValid;
sGtwiz9CtrlAxiBReady <= sGtwiz9CtrlAxiBReady;
sGtwiz9CtrlAxiARAddr <= sGtwiz9CtrlAxiARAddr;
sGtwiz9CtrlAxiARValid <= sGtwiz9CtrlAxiARValid;
sGtwiz9CtrlAxiARReady <= sGtwiz9CtrlAxiARReady;
sGtwiz9CtrlAxiRData <= sGtwiz9CtrlAxiRData;
sGtwiz9CtrlAxiRResp <= sGtwiz9CtrlAxiRResp;
sGtwiz9CtrlAxiRValid <= sGtwiz9CtrlAxiRValid;
sGtwiz9CtrlAxiRReady <= sGtwiz9CtrlAxiRReady;
sGtwiz9DrpChAxiAWAddr <= sGtwiz9DrpChAxiAWAddr;
sGtwiz9DrpChAxiAWValid <= sGtwiz9DrpChAxiAWValid;
sGtwiz9DrpChAxiAWReady <= sGtwiz9DrpChAxiAWReady;
sGtwiz9DrpChAxiWData <= sGtwiz9DrpChAxiWData;
sGtwiz9DrpChAxiWStrb <= sGtwiz9DrpChAxiWStrb;
sGtwiz9DrpChAxiWValid <= sGtwiz9DrpChAxiWValid;
sGtwiz9DrpChAxiWReady <= sGtwiz9DrpChAxiWReady;
sGtwiz9DrpChAxiBResp <= sGtwiz9DrpChAxiBResp;
sGtwiz9DrpChAxiBValid <= sGtwiz9DrpChAxiBValid;
sGtwiz9DrpChAxiBReady <= sGtwiz9DrpChAxiBReady;
sGtwiz9DrpChAxiARAddr <= sGtwiz9DrpChAxiARAddr;
sGtwiz9DrpChAxiARValid <= sGtwiz9DrpChAxiARValid;
sGtwiz9DrpChAxiARReady <= sGtwiz9DrpChAxiARReady;
sGtwiz9DrpChAxiRData <= sGtwiz9DrpChAxiRData;
sGtwiz9DrpChAxiRResp <= sGtwiz9DrpChAxiRResp;
sGtwiz9DrpChAxiRValid <= sGtwiz9DrpChAxiRValid;
sGtwiz9DrpChAxiRReady <= sGtwiz9DrpChAxiRReady;
UserClkPort10 <= UserClkPort10;
aPort10PmaInit <= aPort10PmaInit;
aPort10ResetPb <= aPort10ResetPb;
uPort10AxiTxTData0 <= uPort10AxiTxTData0;
uPort10AxiTxTData1 <= uPort10AxiTxTData1;
uPort10AxiTxTData2 <= uPort10AxiTxTData2;
uPort10AxiTxTData3 <= uPort10AxiTxTData3;
uPort10AxiTxTKeep <= uPort10AxiTxTKeep;
uPort10AxiTxTLast <= uPort10AxiTxTLast;
uPort10AxiTxTValid <= uPort10AxiTxTValid;
uPort10AxiTxTReady <= uPort10AxiTxTReady;
uPort10AxiRxTData0 <= uPort10AxiRxTData0;
uPort10AxiRxTData1 <= uPort10AxiRxTData1;
uPort10AxiRxTData2 <= uPort10AxiRxTData2;
uPort10AxiRxTData3 <= uPort10AxiRxTData3;
uPort10AxiRxTKeep <= uPort10AxiRxTKeep;
uPort10AxiRxTLast <= uPort10AxiRxTLast;
uPort10AxiRxTValid <= uPort10AxiRxTValid;
uPort10AxiNfcTValid <= uPort10AxiNfcTValid;
uPort10AxiNfcTData <= uPort10AxiNfcTData;
uPort10AxiNfcTReady <= uPort10AxiNfcTReady;
uPort10HardError <= uPort10HardError;
uPort10SoftError <= uPort10SoftError;
uPort10LaneUp <= uPort10LaneUp;
uPort10ChannelUp <= uPort10ChannelUp;
uPort10SysResetOut <= uPort10SysResetOut;
uPort10MmcmNotLockOut <= uPort10MmcmNotLockOut;
uPort10CrcPassFail_n <= uPort10CrcPassFail_n;
uPort10CrcValid <= uPort10CrcValid;
iPort10LinkResetOut <= iPort10LinkResetOut;
sGtwiz10CtrlAxiAWAddr <= sGtwiz10CtrlAxiAWAddr;
sGtwiz10CtrlAxiAWValid <= sGtwiz10CtrlAxiAWValid;
sGtwiz10CtrlAxiAWReady <= sGtwiz10CtrlAxiAWReady;
sGtwiz10CtrlAxiWData <= sGtwiz10CtrlAxiWData;
sGtwiz10CtrlAxiWStrb <= sGtwiz10CtrlAxiWStrb;
sGtwiz10CtrlAxiWValid <= sGtwiz10CtrlAxiWValid;
sGtwiz10CtrlAxiWReady <= sGtwiz10CtrlAxiWReady;
sGtwiz10CtrlAxiBResp <= sGtwiz10CtrlAxiBResp;
sGtwiz10CtrlAxiBValid <= sGtwiz10CtrlAxiBValid;
sGtwiz10CtrlAxiBReady <= sGtwiz10CtrlAxiBReady;
sGtwiz10CtrlAxiARAddr <= sGtwiz10CtrlAxiARAddr;
sGtwiz10CtrlAxiARValid <= sGtwiz10CtrlAxiARValid;
sGtwiz10CtrlAxiARReady <= sGtwiz10CtrlAxiARReady;
sGtwiz10CtrlAxiRData <= sGtwiz10CtrlAxiRData;
sGtwiz10CtrlAxiRResp <= sGtwiz10CtrlAxiRResp;
sGtwiz10CtrlAxiRValid <= sGtwiz10CtrlAxiRValid;
sGtwiz10CtrlAxiRReady <= sGtwiz10CtrlAxiRReady;
sGtwiz10DrpChAxiAWAddr <= sGtwiz10DrpChAxiAWAddr;
sGtwiz10DrpChAxiAWValid <= sGtwiz10DrpChAxiAWValid;
sGtwiz10DrpChAxiAWReady <= sGtwiz10DrpChAxiAWReady;
sGtwiz10DrpChAxiWData <= sGtwiz10DrpChAxiWData;
sGtwiz10DrpChAxiWStrb <= sGtwiz10DrpChAxiWStrb;
sGtwiz10DrpChAxiWValid <= sGtwiz10DrpChAxiWValid;
sGtwiz10DrpChAxiWReady <= sGtwiz10DrpChAxiWReady;
sGtwiz10DrpChAxiBResp <= sGtwiz10DrpChAxiBResp;
sGtwiz10DrpChAxiBValid <= sGtwiz10DrpChAxiBValid;
sGtwiz10DrpChAxiBReady <= sGtwiz10DrpChAxiBReady;
sGtwiz10DrpChAxiARAddr <= sGtwiz10DrpChAxiARAddr;
sGtwiz10DrpChAxiARValid <= sGtwiz10DrpChAxiARValid;
sGtwiz10DrpChAxiARReady <= sGtwiz10DrpChAxiARReady;
sGtwiz10DrpChAxiRData <= sGtwiz10DrpChAxiRData;
sGtwiz10DrpChAxiRResp <= sGtwiz10DrpChAxiRResp;
sGtwiz10DrpChAxiRValid <= sGtwiz10DrpChAxiRValid;
sGtwiz10DrpChAxiRReady <= sGtwiz10DrpChAxiRReady;
UserClkPort11 <= UserClkPort11;
aPort11PmaInit <= aPort11PmaInit;
aPort11ResetPb <= aPort11ResetPb;
uPort11AxiTxTData0 <= uPort11AxiTxTData0;
uPort11AxiTxTData1 <= uPort11AxiTxTData1;
uPort11AxiTxTData2 <= uPort11AxiTxTData2;
uPort11AxiTxTData3 <= uPort11AxiTxTData3;
uPort11AxiTxTKeep <= uPort11AxiTxTKeep;
uPort11AxiTxTLast <= uPort11AxiTxTLast;
uPort11AxiTxTValid <= uPort11AxiTxTValid;
uPort11AxiTxTReady <= uPort11AxiTxTReady;
uPort11AxiRxTData0 <= uPort11AxiRxTData0;
uPort11AxiRxTData1 <= uPort11AxiRxTData1;
uPort11AxiRxTData2 <= uPort11AxiRxTData2;
uPort11AxiRxTData3 <= uPort11AxiRxTData3;
uPort11AxiRxTKeep <= uPort11AxiRxTKeep;
uPort11AxiRxTLast <= uPort11AxiRxTLast;
uPort11AxiRxTValid <= uPort11AxiRxTValid;
uPort11AxiNfcTValid <= uPort11AxiNfcTValid;
uPort11AxiNfcTData <= uPort11AxiNfcTData;
uPort11AxiNfcTReady <= uPort11AxiNfcTReady;
uPort11HardError <= uPort11HardError;
uPort11SoftError <= uPort11SoftError;
uPort11LaneUp <= uPort11LaneUp;
uPort11ChannelUp <= uPort11ChannelUp;
uPort11SysResetOut <= uPort11SysResetOut;
uPort11MmcmNotLockOut <= uPort11MmcmNotLockOut;
uPort11CrcPassFail_n <= uPort11CrcPassFail_n;
uPort11CrcValid <= uPort11CrcValid;
iPort11LinkResetOut <= iPort11LinkResetOut;
sGtwiz11CtrlAxiAWAddr <= sGtwiz11CtrlAxiAWAddr;
sGtwiz11CtrlAxiAWValid <= sGtwiz11CtrlAxiAWValid;
sGtwiz11CtrlAxiAWReady <= sGtwiz11CtrlAxiAWReady;
sGtwiz11CtrlAxiWData <= sGtwiz11CtrlAxiWData;
sGtwiz11CtrlAxiWStrb <= sGtwiz11CtrlAxiWStrb;
sGtwiz11CtrlAxiWValid <= sGtwiz11CtrlAxiWValid;
sGtwiz11CtrlAxiWReady <= sGtwiz11CtrlAxiWReady;
sGtwiz11CtrlAxiBResp <= sGtwiz11CtrlAxiBResp;
sGtwiz11CtrlAxiBValid <= sGtwiz11CtrlAxiBValid;
sGtwiz11CtrlAxiBReady <= sGtwiz11CtrlAxiBReady;
sGtwiz11CtrlAxiARAddr <= sGtwiz11CtrlAxiARAddr;
sGtwiz11CtrlAxiARValid <= sGtwiz11CtrlAxiARValid;
sGtwiz11CtrlAxiARReady <= sGtwiz11CtrlAxiARReady;
sGtwiz11CtrlAxiRData <= sGtwiz11CtrlAxiRData;
sGtwiz11CtrlAxiRResp <= sGtwiz11CtrlAxiRResp;
sGtwiz11CtrlAxiRValid <= sGtwiz11CtrlAxiRValid;
sGtwiz11CtrlAxiRReady <= sGtwiz11CtrlAxiRReady;
sGtwiz11DrpChAxiAWAddr <= sGtwiz11DrpChAxiAWAddr;
sGtwiz11DrpChAxiAWValid <= sGtwiz11DrpChAxiAWValid;
sGtwiz11DrpChAxiAWReady <= sGtwiz11DrpChAxiAWReady;
sGtwiz11DrpChAxiWData <= sGtwiz11DrpChAxiWData;
sGtwiz11DrpChAxiWStrb <= sGtwiz11DrpChAxiWStrb;
sGtwiz11DrpChAxiWValid <= sGtwiz11DrpChAxiWValid;
sGtwiz11DrpChAxiWReady <= sGtwiz11DrpChAxiWReady;
sGtwiz11DrpChAxiBResp <= sGtwiz11DrpChAxiBResp;
sGtwiz11DrpChAxiBValid <= sGtwiz11DrpChAxiBValid;
sGtwiz11DrpChAxiBReady <= sGtwiz11DrpChAxiBReady;
sGtwiz11DrpChAxiARAddr <= sGtwiz11DrpChAxiARAddr;
sGtwiz11DrpChAxiARValid <= sGtwiz11DrpChAxiARValid;
sGtwiz11DrpChAxiARReady <= sGtwiz11DrpChAxiARReady;
sGtwiz11DrpChAxiRData <= sGtwiz11DrpChAxiRData;
sGtwiz11DrpChAxiRResp <= sGtwiz11DrpChAxiRResp;
sGtwiz11DrpChAxiRValid <= sGtwiz11DrpChAxiRValid;
sGtwiz11DrpChAxiRReady <= sGtwiz11DrpChAxiRReady;