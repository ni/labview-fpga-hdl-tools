-------------------------------------------------------------------------------
--
-- File: PkgLvFpgaConst.vhd
-- Author: David Cabrera
-- Original Project: Puma K7
-- Date: 22 July 2013
--
-------------------------------------------------------------------------------
-- (c) 2025 Copyright National Instruments Corporation
-- 
-- SPDX-License-Identifier: MIT
-------------------------------------------------------------------------------
--
-- Purpose:
--  This file will be generated by LV FPGA to set constants required for
--  Puma K7 compilation.
--
-------------------------------------------------------------------------------
--
-- githubvisible=true

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package PkgLvFpgaConst is

  -----------------------------------------------------------------------------
  -- LV FPGA generated constants
  -----------------------------------------------------------------------------

  constant kExpectedTbId   : std_logic_vector(31 downto 0) := X"D00FD00F";
  constant kExpectDumbTb   : std_logic := '1';
  constant kEnableFamClockSync : std_logic := '0';
  constant kFamClockSrcSel  : std_logic := '0';
  constant kInsertBank0Mig  : boolean := false;
  constant kInsertBank1Mig  : boolean := false;
  constant kAuxDioDefaultVoltage : natural := 3300;
  constant kAuxMgtClipPresent : boolean := false;
  constant kCfgSubsysId : std_logic_vector(15 downto 0) := X"78F9";  

  -- Required for HMB
  constant kDram2DPBaseAddress : natural := 16#20000#;
  constant kInsertHostMemoryBufferMig : boolean := false;
  constant kInsertLowLatencyBufferMig : boolean := false;

end PkgLvFpgaConst;

package body PkgLvFpgaConst is

  
end PkgLvFpgaConst;

